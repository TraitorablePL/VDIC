package shape_pkg;

`include "shape.svh"
`include "rectangle.svh"
`include "square.svh"
`include "triangle.svh"
`include "shape_factory.svh"
`include "shape_reporter.svh"

endpackage : shape_pkg