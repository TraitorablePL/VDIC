class Extreme_val_command extends Random_command;
    
    `uvm_object_utils(Extreme_val_command)
    

// Constraints

    //TODO
        
// Command transaction constructor
 
    function new(string name = "");
        super.new(name);
    endfunction : new
    
endclass : Extreme_val_command